module and_gate (
    input logic zero_flag,      
    input logic branch,      
    output logic PCsrc 
);

    assign result = a & b;  // Bitwise AND operation

endmodule
